otutay@eotPc.18126:1615923773