package packageTb;
   localparam logic [5:0]  Rtype = 6'b000001;
   localparam logic [5:0]  Itype = 6'b000010;
   localparam logic [5:0]  Stype = 6'b000100;
   localparam logic [5:0]  Btype = 6'b001000;
   localparam logic [5:0]  Utype = 6'b010000;
   localparam logic [5:0]  Jtype = 6'b100000;




endpackage : packageTb
