-------------------------------------------------------------------------------
-- Title      : fetchWB
-- Project    :
-------------------------------------------------------------------------------
-- File       : fetchWb.vhd
-- Author     : osmant  <otutaysalgir@gmail.com>
-- Company    :
-- Created    : 2021-03-25
-- Last update: 2021-03-26
-- Platform   :
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: fetch wb stage
-------------------------------------------------------------------------------
-- Copyright (c) 2021
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2021-03-25  1.0      otutay	Created
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.corePckg.all;

entity fetchWb is

  port (
    iClk : in std_logic
    );

end entity fetchWb;

architecture rtl of fetchWb is

begin  -- architecture rtl



end architecture rtl;
