otutay@eotPc.2502:1615923773